`default_nettype none     // Disable implicit nets. Reduces some types of bugs.
module top_module( 
    input wire [15:0] in,
    output wire [7:0] out_hi,
    output wire [7:0] out_lo );
    // Split the 16-bit input into two 8-bit outputs using concatenation
    assign {out_hi, out_lo} = in;

    // Alternative approach using explicit bit slicing:
    // assign out_hi = in[15:8];
    // assign out_lo = in[7:0];
endmodule
